Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

Entity Time_RUN is
End Time_RUN;

architecture Behavioral of Time_RUN is

begin


end Behavioral;

